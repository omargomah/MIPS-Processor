
library ieee;
use ieee.std_logic_1164.all;
entity Mux is
    port (
       A: in  std_logic_vector(31 downto 0);
       B: in  std_logic_vector(31 downto 0);
       Sel: in  std_logic;
       Y: out std_logic_vector(31 downto 0));
end  Mux ;
architecture behavier of Mux  is
begin
    Y<= B when Sel = '1' else A;
end behavier;
