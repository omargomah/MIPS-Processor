library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity Adder is
    port (  
        A: in  std_logic_vector(31 downto 0);
        B: in  std_logic_vector(31 downto 0);
       Sum: out std_logic_vector(31 downto 0));
end entity Adder;
architecture Behavioral of Adder is
begin
    Sum <= std_logic_vector(signed(A) + signed(B));
end architecture Behavioral;
